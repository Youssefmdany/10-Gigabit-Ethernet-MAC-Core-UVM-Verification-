

class Base_Sequence extends uvm_sequence #(Packet);




   `uvm_object_utils(Base_Sequence)
	
	

	
	
	
	
	function new (string name = "Base_Sequence");
	
	
	    super.new(name); 
	
	
	endfunction: new

	
	
	
	


endclass: Base_Sequence